module dec_2x4(y,a,b,en); 
    input a,b,en; 
    output reg [3:0]y; 

    always @(a,b,en)
        begin
            if (en==0)
                begin
                    if(a==1'b0 & b==1'b0) 
                        y=4'b1110; 
                    else if(a==1'b0 & b==1'b1) 
                        y=4'b1101; 
                    else if(a==1'b1 & b==1'b0) 
                        y=4'b1011; 
                    else if(a==1'b1 & b==1'b1) 
                        y=4'b0111; 
                    else 
                        y=4'bxxxx;
                end
            else 
                y=4'b1111;
        end
endmodule